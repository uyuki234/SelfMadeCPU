module adder8_tb;
    reg             clk = 1'b0;
    reg     [7:0]   in0 = 8'h00;
    reg     [7:0]   in1 = 8'h00;
    wire    [7:0]   out;

    initial begin
        $dumpfile("wave.vcd");
        $dumpvars(0, DUT);
    end

    always #1 begin
        clk <= ~clk;
    end

    adder8 DUT(
        .clk    (clk    ),
        .in0    (in0    ),
        .in1    (in1    ),
        .out    (out    )
    );

    initial begin
        #2
        in0 = 8'h05;
        in1 = 8'h04;
        #2
        in0 = 8'hff;
        in1 = 8'h01;
        #2
        $finish;
    end
endmodule
